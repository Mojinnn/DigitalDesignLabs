library verilog;
use verilog.vl_types.all;
entity CodeVHDL_vlg_vec_tst is
end CodeVHDL_vlg_vec_tst;
