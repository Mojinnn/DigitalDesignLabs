library verilog;
use verilog.vl_types.all;
entity CongOR_vlg_vec_tst is
end CongOR_vlg_vec_tst;
