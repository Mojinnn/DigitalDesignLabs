library verilog;
use verilog.vl_types.all;
entity CongNOT_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CongNOT_vlg_check_tst;
