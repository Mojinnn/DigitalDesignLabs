library verilog;
use verilog.vl_types.all;
entity CongNOT_vlg_vec_tst is
end CongNOT_vlg_vec_tst;
