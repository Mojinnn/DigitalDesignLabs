library verilog;
use verilog.vl_types.all;
entity KTS_vlg_check_tst is
    port(
        O               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end KTS_vlg_check_tst;
