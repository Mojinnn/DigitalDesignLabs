library verilog;
use verilog.vl_types.all;
entity CongAND_vlg_check_tst is
    port(
        O               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CongAND_vlg_check_tst;
