library verilog;
use verilog.vl_types.all;
entity CongAND_vlg_vec_tst is
end CongAND_vlg_vec_tst;
