library verilog;
use verilog.vl_types.all;
entity KTS_vlg_vec_tst is
end KTS_vlg_vec_tst;
